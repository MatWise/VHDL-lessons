architecture behav of analyzer is
begin
  process is
    variable cycle_length_counter: integer;
    variable start_value: std_logic_vector(7 downto 0);
  begin
    wait until res_n = '1';
    loop
      wait on clk until clk = '1' and reset = '1';
      cycle_length_counter := 1;
      wait on clk until clk = '1' and reset = '0';
      start_value := q;
      wait on clk until clk = '1';
      while q /= start_value loop
        cycle_length_counter := cycle_length_counter + 1;
        wait on clk until clk = '1';
      end loop;
      report "cycle length: " & integer'image(cycle_length_counter);
    end loop;
  end process;
end architecture behav; 