library ieee; use ieee.std_logic_1164.all;

entity galois_analyzer is
  port(
    clk: in std_logic;
    res_n: in std_logic;
    reset: in std_logic;
    q: in std_logic_vector(7 downto 0));
end entity galois_analyzer;
