entity galois_lfsr_tb is
end entity galois_lfsr_tb;
