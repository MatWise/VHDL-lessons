entity senso is
end entity senso;
