entity random_tb is
end entity random_tb;
