architecture behav of timer is
begin
  process(clk, res_n) is
    

end architecture behav;