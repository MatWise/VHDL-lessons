entity timer_tb is
end entity timer_tb;
