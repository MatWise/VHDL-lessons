entity counter_tb is
end entity counter_tb;
