entity button_tb is
end entity button_tb;
