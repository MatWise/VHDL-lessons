library ieee; use ieee.std_logic_1164.all;

entity clk_res_gen is
  port(
    clk, res_n: out std_logic);
end entity clk_res_gen;
