library ieee; use ieee.std_logic_1164.all;

entity button_tester is
  port(
    tx_n: out std_logic);
end entity button_tester;
